.include '45nm_LP.pm'

.SUBCKT PC BL BLB PRE Vdd
M_i_2 BL PRE Vvdd Vdd PMOS_VTL W=0.630000U L=0.050000U
M_i_3 BLB PRE Vvdd Vdd PMOS_VTL W=0.630000U L=0.050000U
M_i_4 BL PRE BLB Vdd PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

