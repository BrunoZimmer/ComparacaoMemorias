*transmission gate

.SUBCKT TG IN ZN EN VDD VSS
*M_i Drain Gate Source Bulk
M_i_2 IN EN ZN VSS NMOS W=15.15000U L=0.050000U

M_i_3 IN ENB ZN VDD PMOS W=30.630000U L=0.050000U

M_i_6 EN ENB VDD VDD PMOS W=4.630000U L=0.050000U
M_i_7 EN ENB VSS VSS NMOS W=8.630000U L=0.050000U
.ENDS 
