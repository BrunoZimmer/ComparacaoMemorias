*.include '45nm_LP.pm'

.SUBCKT INV A ZN VDD VSS 
*M_i Drain Gate Source Bulk
M_i_0 ZN A VSS VSS NMOS_VTL W=0.415000U L=0.050000U
M_i_1 ZN A VDD VDD PMOS_VTL W=0.630000U L=0.050000U
.ENDS 

