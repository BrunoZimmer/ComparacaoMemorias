*tristate
.include 'MTJT.spi'

.SUBCKT BCTM BL SL WL
X1 NM BL MTJT
M_i_1 NM WL SL SL PMOS W=12.630000U L=0.050000U
.ENDS 

